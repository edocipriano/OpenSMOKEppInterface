   THERMO 
   300.0   1000.0   3000.0
N2                G 8/02N   2    0    0    0G   200.000  6000.00  1000.00      1
 2.95257637E+00 1.39690040E-03-4.92631603E-07 7.86010195E-11-4.60755204E-15    2
-9.23948688E+02 5.87188762E+00 3.53100528E+00-1.23660988E-04-5.02999433E-07    3
 2.43530612E-09-1.40881235E-12-1.04697628E+03 2.96747038E+00 0.00000000E+00    4
P-HDPE-P                C  40H  80          G    200.00   2000.00 1500.00      1
 9.46552181E+01 1.48843812E-01 8.28388378E-05-9.89931381E-08 2.32390625E-11    2
-1.60002354E+05-4.14345049E+02 9.46552181E+01 1.48843812E-01 8.28388378E-05    3
-9.89931381E-08 2.32390625E-11-1.60002354E+05-4.14345049E+02                   4
C2H4                    C   2H   4          G    300.00   4000.00 1000.00      1
 .399182724E+01 .104833908E-01-.371721342E-05 .594628366E-09-.353630386E-13    2
 .426865851E+04-.269081762E+00 .395920063E+01-.757051373E-02 .570989993E-04    3
-.691588352E-07 .269884190E-10 .508977598E+04 .409730213E+01                   4
