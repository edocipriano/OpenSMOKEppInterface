! This thermodynamic database was obtained by fitting the thermodynamic properties
! extracted from the following file: CRECK_2003_C1_C3_HT.CKT
! The thermodynamic properties are fitted in order to preserve not only the 
! continuity of each function at the intermediate temperature, but also the  continuity
! of the derivatives, from the 1st to the 3rd order
! The intermediate temperatures are the same for all the species.
! Last update: 11/26/2023

THERMO ALL
270.   1000.   3500. 
CH3OH                   C   1H   4O   1     G    300.00   3500.00 1000.00      1
 1.36199082e+00 1.47016350e-02-6.74192919e-06 1.50725057e-09-1.33717354e-13    2
-2.52166926e+04 1.70048495e+01 6.28410461e-01 1.76359564e-02-1.11434113e-05    3
 4.44157201e-09-8.67297713e-13-2.50699765e+04 2.05439507e+01                   4
H2                      H   2               G    200.00   3500.00 1000.00      1
 4.06077528e+00-1.67367616e-03 1.75993108e-06-5.86430223e-10 6.65899071e-14    2
-1.18864369e+03-7.08382230e+00 2.98310117e+00 2.63702026e-03-4.70611354e-06    3
 3.72426619e-09-1.01108420e-12-9.73108868e+02-1.88466771e+00                   4
H                       H   1               G    200.00   3500.00 1000.00      1
 2.50043469e+00-1.05089320e-06 8.56597149e-10-2.82344590e-13 3.23453433e-17    2
 2.54736098e+04-4.48994333e-01 2.49958759e+00 2.33750216e-06-4.22599589e-09    3
 3.10605077e-12-8.14753497e-16 2.54737793e+04-4.44907570e-01                   4
O2                      O   2               G    200.00   3500.00 1000.00      1
 2.59418011e+00 3.01293505e-03-1.93158331e-06 5.84246115e-10-6.41585618e-14    2
-8.61799675e+02 9.14749788e+00 3.46761808e+00-4.80816814e-04 3.30904448e-06    3
-2.90950575e-09 8.09279404e-13-1.03648727e+03 4.93366459e+00                   4
O                       O   1               G    200.00   3500.00 1000.00      1
 2.50077543e+00 8.39962383e-05-9.75880148e-08 3.62707395e-11-4.12114418e-15    2
 2.92445463e+04 5.14506503e+00 3.00716588e+00-1.94156558e-03 2.94075471e-06    3
-1.98929107e-09 5.02269309e-13 2.91432682e+04 2.70202381e+00                   4
H2O                     H   2O   1          G    200.00   3500.00 1000.00      1
 3.30588708e+00 1.74342157e-03 5.12337364e-08-1.46310042e-10 2.14519038e-14    2
-3.01205579e+04 3.43022225e+00 4.17881168e+00-1.74827683e-03 5.28878133e-06    3
-3.63800844e-09 8.94376503e-13-3.02951428e+04-7.81134343e-01                   4
OH                      H   1O   1          G    200.00   3500.00 1000.00      1
 3.47656309e+00-2.30512504e-04 6.85003016e-07-2.58084516e-10 3.04253084e-14    2
 3.49661263e+03 2.38083066e+00 4.00594686e+00-2.34804762e-03 3.86130568e-06    3
-2.37561963e-09 5.59809087e-13 3.39073587e+03-1.73140053e-01                   4
H2O2                    H   2O   2          G    200.00   3500.00 1000.00      1
 3.69620772e+00 5.92424119e-03-2.59473223e-06 5.93112571e-10-5.42682448e-14    2
-1.76560131e+04 5.44017070e+00 3.26921550e+00 7.63221008e-03-5.15668557e-06    3
 2.30108146e-09-4.81260468e-13-1.75706147e+04 7.50016135e+00                   4
HO2                     H   1O   2          G    200.00   3500.00 1000.00      1
 2.87816085e+00 4.80634573e-03-2.50212755e-06 7.00245313e-10-7.63793313e-14    2
 4.44209110e+02 9.88006528e+00 3.44162180e+00 2.55250194e-03 8.78638140e-07    3
-1.55359848e-09 4.87081617e-13 3.31516920e+02 7.16169191e+00                   4
CO                      C   1O   1          G    200.00   3500.00 1000.00      1
 2.74907495e+00 1.97367768e-03-9.36103965e-07 2.15530966e-10-1.95219158e-14    2
-1.41583305e+04 7.64673793e+00 3.73475699e+00-1.96905047e-03 4.97798827e-06    3
-3.72719719e-09 9.66160123e-13-1.43554669e+04 2.89139187e+00                   4
CO2                     C   1O   2          G    200.00   3500.00 1000.00      1
 3.54460780e+00 5.01221005e-03-2.64865077e-06 6.65160387e-10-6.42432119e-14    2
-4.86279535e+04 4.01016765e+00 2.11557108e+00 1.07283569e-02-1.12228711e-05    3
 6.38130728e-09-1.49327994e-12-4.83421461e+04 1.09044438e+01                   4
CH4                     C   1H   4          G    300.00   3500.00 1000.00      1
-1.03344835e-01 1.37591208e-02-6.07522307e-06 1.38758156e-09-1.24974791e-13    2
-9.39493046e+03 1.94243232e+01 2.95013182e+00 1.54521422e-03 1.22456369e-05    3
-1.08263251e-08 2.92850187e-12-1.00056258e+04 4.69306337e+00                   4
CH3                     C   1H   3          G    300.00   3500.00 1000.00      1
 2.82634627e+00 6.06830643e-03-2.14837164e-06 3.54546043e-10-2.26100123e-14    2
 1.65733843e+04 5.57284900e+00 3.51500165e+00 3.31368488e-03 1.98356069e-06    3
-2.40007551e-09 6.66045375e-13 1.64356532e+04 2.25048484e+00                   4
CH2                     C   1H   2          G    300.00   3500.00 1000.00      1
 3.50279627e+00 2.25680851e-03-4.11311887e-07-3.16119544e-11 1.15424126e-14    2
 4.59259048e+04 2.80775303e+00 3.87638279e+00 7.62462421e-04 1.83020725e-06    3
-1.52595804e-09 3.85128935e-13 4.58511875e+04 1.00541401e+00                   4
CH2(S)                  C   1H   2          G    300.00   3500.00 1000.00      1
 2.72267961e+00 3.73668496e-03-1.41857410e-06 2.94773602e-10-2.58912481e-14    2
 5.06549560e+04 6.31301629e+00 4.13684563e+00-1.91997915e-03 7.06642206e-06    3
-5.36189051e-09 1.38827478e-12 5.03721228e+04-5.09517328e-01                   4
CH3O                    C   1H   3O   1     G    300.00   3500.00 1000.00      1
 2.41318476e+00 1.22101388e-02-6.11028600e-06 1.46676389e-09-1.37436418e-13    2
 1.24867034e+03 1.08490945e+01 2.65211891e-01 2.08020303e-02-1.89981232e-05    3
 1.00586554e-08-2.28540929e-12 1.67826492e+03 2.12118220e+01                   4
CH2OH                   C   1H   3O   1     G    300.00   3500.00 1000.00      1
 4.08435451e+00 8.00757963e-03-3.54698535e-06 7.71850004e-10-6.74865850e-14    2
-3.68580525e+03 3.66682075e+00 1.89045633e+00 1.67831723e-02-1.67103744e-05    3
 9.54744271e-09-2.26138476e-12-3.24702562e+03 1.42511113e+01                   4
CH2O                    C   1H   2O   1     G    300.00   3500.00 1000.00      1
 9.48565662e-01 1.09688025e-02-5.81045395e-06 1.47149667e-09-1.44094288e-13    2
-1.37848123e+04 1.80455343e+01 2.87885429e+00 3.24764803e-03 5.77127783e-06    3
-6.24965785e-09 1.78619434e-12-1.41708700e+04 8.73300751e+00                   4
HCO                     C   1H   1O   1     G    200.00   3500.00 1000.00      1
 2.29086776e+00 6.01826018e-03-3.26408994e-06 9.06148666e-10-9.53398930e-14    2
 4.15288903e+03 1.23882062e+01 3.74614032e+00 1.97169955e-04 5.46754540e-06    3
-4.91494156e-09 1.35993266e-12 3.86183452e+03 5.36735734e+00                   4
C2H4                    C   2H   4          G    300.00   3500.00 1000.00      1
 1.72159882e+00 1.51093228e-02-7.03615661e-06 1.59719862e-09-1.43847181e-13    2
 5.10084649e+03 1.21382035e+01-7.43812044e-01 2.49709662e-02-2.18286218e-05    3
 1.14588421e-08-2.60925805e-12 5.59392866e+03 2.40323857e+01                   4
C2H3                    C   2H   3          G    300.00   3500.00 1000.00      1
 2.87744740e+00 1.01276366e-02-4.48501948e-06 9.76327127e-10-8.51883496e-14    2
 3.43280675e+04 8.69075318e+00 7.28453850e-01 1.87236108e-02-1.73789808e-05    3
 9.57230133e-09-2.23418190e-12 3.47578663e+04 1.90584048e+01                   4
N2                      N   2               G    200.00   3500.00 1000.00      1
 2.86445153e+00 1.55307425e-03-5.90242371e-07 1.04543577e-10-7.10938713e-15    2
-8.87270169e+02 6.36509032e+00 3.75301206e+00-2.00116785e-03 4.74112078e-06    3
-3.44969853e-09 8.81451139e-13-1.06498227e+03 2.07829942e+00                   4
END
