! This thermodynamic database was obtained by fitting the thermodynamic properties
! extracted from the following file: CRECK_2003_C1_C3_HT.CKT
! The thermodynamic properties are fitted in order to preserve not only the 
! continuity of each function at the intermediate temperature, but also the  continuity
! of the derivatives, from the 1st to the 3rd order
! The intermediate temperatures are chosen in order to minimize the fitting error.
! Last update: 11/26/2023

THERMO ALL
270.   1000.   3500. 
CH3OH                   C   1H   4O   1     G    300.00   3500.00 1800.00      1
 2.71701641e+00 1.21538330e-02-5.02106867e-06 1.01068022e-09-8.18460330e-14    2
-2.57693414e+04 9.47419935e+00 8.47330413e-01 1.63086907e-02-8.48345015e-06    3
 2.29304373e-09-2.59952076e-13-2.50962544e+04 1.95933300e+01                   4
H2                      H   2               G    200.00   3500.00  700.00      1
 3.78199882e+00-1.01873266e-03 1.24226241e-06-4.19011929e-10 4.75543833e-14    2
-1.10283023e+03-5.60525911e+00 2.64204442e+00 5.49529249e-03-1.27163629e-05    3
 1.28749170e-08-4.70027736e-12-9.43236618e+02-5.12231254e-01                   4
H                       H   1               G    200.00   3500.00  860.00      1
 2.50031492e+00-7.73402937e-07 6.39349536e-10-2.12554688e-13 2.44483709e-17    2
 2.54736474e+04-4.48357209e-01 2.49950545e+00 2.99160533e-06-5.92752534e-09    3
 4.87804599e-12-1.45537741e-15 2.54737866e+04-4.44574039e-01                   4
O2                      O   2               G    200.00   3500.00  700.00      1
 2.82012408e+00 2.48211357e-03-1.51202094e-06 4.48556199e-10-4.87305665e-14    2
-9.31350152e+02 7.94914552e+00 3.74403921e+00-2.79740146e-03 9.80122556e-06    3
-1.03259643e-08 3.79931246e-12-1.06069827e+03 3.82132646e+00                   4
O                       O   1               G    200.00   3500.00  720.00      1
 2.62549143e+00-2.08959638e-04 1.33918542e-07-3.85875887e-11 4.38918680e-15    2
 2.92061519e+04 4.48358521e+00 3.14799201e+00-3.11174067e-03 6.18137903e-06    3
-5.63808804e-09 1.94866018e-12 2.91309118e+04 2.13446548e+00                   4
H2O                     H   2O   1          G    200.00   3500.00 1420.00      1
 2.66777069e+00 3.05768864e-03-9.00442530e-07 1.43361590e-10-1.00857860e-14    2
-2.98875645e+04 6.91191161e+00 4.06061173e+00-8.65807224e-04 3.24409535e-06    3
-1.80243084e-09 3.32483304e-13-3.02831314e+04-2.96150501e-01                   4
OH                      H   1O   1          G    200.00   3500.00 1700.00      1
 2.49867381e+00 1.66635254e-03-6.28251336e-07 1.28346754e-10-1.05735839e-14    2
 3.88110712e+03 7.78218797e+00 3.91354630e+00-1.66275921e-03 2.30920021e-06    3
-1.02359503e-09 1.58829619e-13 3.40005047e+03 2.05474752e-01                   4
H2O2                    H   2O   2          G    200.00   3500.00 1800.00      1
 4.76869611e+00 3.89237905e-03-1.21382388e-06 1.92615393e-10-1.22582099e-14    2
-1.80900219e+04-5.11810218e-01 3.34774226e+00 7.05005427e-03-3.84521989e-06    3
 1.16720651e-09-1.47618087e-13-1.75784785e+04 7.17868844e+00                   4
HO2                     H   1O   2          G    200.00   3500.00  700.00      1
 3.02391888e+00 4.46390907e-03-2.23146491e-06 6.12710795e-10-6.64266231e-14    2
 3.99341609e+02 9.10699973e+00 3.61994300e+00 1.05805700e-03 5.06678953e-06    3
-6.33800772e-09 2.41597285e-12 3.15898233e+02 6.44411479e+00                   4
CO                      C   1O   1          G    200.00   3500.00  960.00      1
 2.79255379e+00 1.87486889e-03-8.59711939e-07 1.91200073e-10-1.67855288e-14    2
-1.41723335e+04 7.41443567e+00 3.75723892e+00-2.14465247e-03 5.42079018e-06    3
-4.17025973e-09 1.11901130e-12-1.43575530e+04 2.79976795e+00                   4
CO2                     C   1O   2          G    200.00   3500.00 1450.00      1
 4.70876459e+00 2.62914723e-03-9.30606600e-07 1.43892961e-10-7.62581846e-15    2
-4.90562638e+04-2.34976404e+00 2.31684348e+00 9.22755029e-03-7.75654080e-06    3
 3.28225351e-09-5.48722465e-13-4.83626067e+04 1.00786234e+01                   4
CH4                     C   1H   4          G    300.00   3500.00  700.00      1
 5.05346503e-01 1.23697842e-02-4.99807899e-06 1.04392757e-09-8.62897323e-14    2
-9.58982505e+03 1.61752770e+01 5.23967302e+00-1.46835102e-02 5.29732662e-05    3
-5.41668773e-08 1.96318549e-11-1.02526308e+04-4.97649608e+00                   4
CH3                     C   1H   3          G    300.00   3500.00 1060.00      1
 2.78805103e+00 6.15233477e-03-2.21179348e-06 3.74402643e-10-2.48151342e-14    2
 1.65862829e+04 5.77899820e+00 3.47829311e+00 3.54764767e-03 1.47408448e-06    3
-1.94375960e-09 5.21921244e-13 1.64399516e+04 2.40875951e+00                   4
CH2                     C   1H   2          G    300.00   3500.00 1800.00      1
 2.81272979e+00 3.55431373e-03-1.28768512e-06 2.21273711e-10-1.48738112e-14    2
 4.62073492e+04 6.64284613e+00 3.76489460e+00 1.43839193e-03 4.75583051e-07    3
-4.31788574e-10 7.58292840e-14 4.58645699e+04 1.48953154e+00                   4
CH2(S)                  C   1H   2          G    300.00   3500.00  970.00      1
 2.75934297e+00 3.65468310e-03-1.35589915e-06 2.74980414e-10-2.36795474e-14    2
 5.06429079e+04 6.11646390e+00 4.18185436e+00-2.21134323e-03 7.71527558e-06    3
-5.95950394e-09 1.58314632e-12 5.03669407e+04-7.03002672e-01                   4
CH3O                    C   1H   3O   1     G    300.00   3500.00 1740.00      1
 5.72238202e+00 5.90227348e-03-1.80340517e-06 2.13334417e-10-5.61810225e-15    2
-7.86257462e+01-7.49174438e+00 8.89660877e-01 1.70119773e-02-1.13807360e-05    3
 3.88280984e-09-5.32841582e-13 1.60316121e+03 1.85001139e+01                   4
CH2OH                   C   1H   3O   1     G    300.00   3500.00 1360.00      1
 5.04534889e+00 6.02727212e-03-2.11386943e-06 3.36086293e-10-2.00987914e-14    2
-4.03584125e+03-1.57523751e+00 2.34821588e+00 1.39600163e-02-1.08632196e-05    3
 4.62498344e-09-8.08499002e-13-3.30222107e+03 1.22661973e+01                   4
CH2O                    C   1H   2O   1     G    300.00   3500.00  700.00      1
 1.33335654e+00 1.00905182e-02-5.12952556e-06 1.25425205e-09-1.19639106e-13    2
-1.39080170e+04 1.59916143e+01 4.32621280e+00-7.01151755e-03 3.15176940e-05    3
-3.36478618e-08 1.23454016e-11-1.43270169e+04 2.62028972e+00                   4
HCO                     C   1H   1O   1     G    200.00   3500.00  770.00      1
 2.60049318e+00 5.29278251e-03-2.69184203e-06 7.21357765e-10-7.43521367e-14    2
 4.05725330e+03 1.07450933e+01 4.03483983e+00-2.15836887e-03 1.18233879e-05    3
-1.18459409e-08 4.00593964e-12 3.83636392e+03 4.20008755e+00                   4
C2H4                    C   2H   4          G    300.00   3500.00 1650.00      1
 4.60402728e+00 9.50595335e-03-3.15129253e-06 4.53052054e-10-2.23949142e-14    2
 3.97229098e+03-3.77420958e+00-6.02932629e-02 2.08133971e-02-1.34307868e-05    3
 4.60638309e-09-6.51687495e-13 5.51151676e+03 2.10642173e+01                   4
C2H3                    C   2H   3          G    300.00   3500.00 1450.00      1
 4.18728253e+00 7.47581889e-03-2.58984461e-06 4.05266527e-10-2.35023527e-14    2
 3.38403788e+04 1.51959400e+00 1.23421229e+00 1.56222195e-02-1.10171556e-05    3
 4.27989229e-09-6.91541277e-13 3.46967692e+04 1.68637042e+01                   4
N2                      N   2               G    200.00   3500.00 1050.00      1
 2.81166073e+00 1.67067353e-03-6.79997421e-07 1.32881376e-10-1.02767438e-14    2
-8.69811581e+02 6.64838048e+00 3.73100682e+00-1.83159730e-03 4.32324661e-06    3
-3.04378150e-09 7.46071560e-13-1.06287426e+03 2.16821198e+00                   4
END
