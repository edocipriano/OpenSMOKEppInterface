   THERMO 
   300.0   1000.0   3000.0
N2                G 8/02N   2    0    0    0G   200.000  6000.00  1000.00      1
 2.95257637E+00 1.39690040E-03-4.92631603E-07 7.86010195E-11-4.60755204E-15    2
-9.23948688E+02 5.87188762E+00 3.53100528E+00-1.23660988E-04-5.02999433E-07    3
 2.43530612E-09-1.40881235E-12-1.04697628E+03 2.96747038E+00 0.00000000E+00    4
BIOMASS                 C   6H  10O   5     S 300.0    4000.0    1000.0        1!From CELL
 2.92516210e+01 1.95010807e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-1.25919988e+05 0.00000000e+00 2.92516210e+01 1.95010807e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-1.25919988e+05 0.00000000e+00                   4
H2O               ATcT3EH   2O   1    0    0G    200.00   6000.00 1000.00      1
 2.73117512E+00 2.95136995E-03-8.35359785E-07 1.26088593E-10-8.40531676E-15    2
-2.99169082E+04 6.55183000E+00 4.20147551E+00-2.05583546E-03 6.56547207E-06    3
-5.52906960E-09 1.78282605E-12-3.02950066E+04-8.60610906E-01-2.90858262E+04    4
CHAR                    C   1               S 300.0    4000.0    1000.0        1
-1.00796361E-01	4.99828606E-03 0.00000000E+00 0.00000000E+00 0.00000000E+00    2           
-1.94683964E+02 0.00000000E+00-1.00796361E-01 4.99828606E-03 0.00000000E+00    3
 0.00000000E+00	0.00000000E+00-1.94683964E+02 0.00000000E+00                   4
TAR                     C   6H  10O   5     S 300.0    4000.0    1000.0        1!From CELL
 .279850422E+02 .264166682E-01-.913640739E-05 .142923991E-08-.833656585E-13    2
-.114313686E+06-.117754445E+03-.781241700E+01 .125424511E+00-.116271866E-03    3
 .544734561E-07-.100746170E-10-.103428291E+06 .690300863E+02                   4

