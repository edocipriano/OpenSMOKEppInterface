! This thermodynamic database was obtained by fitting the thermodynamic properties
! extracted from the following file: CRECK_2003_C1_C3_HT.CKT
! The thermodynamic properties are fitted in order to preserve not only the 
! continuity of each function at the intermediate temperature, but also the  continuity
! of the derivatives, from the 1st to the 3rd order
! The intermediate temperatures are chosen in order to minimize the fitting error.
! Last update: 12/4/2023

THERMO ALL
270.   1000.   3500. 
C2H5OH                  C   2H   6O   1     G    300.00   3500.00 1580.00      1
 7.32490782e+00 1.39762986e-02-4.67366813e-06 6.82063871e-10-3.47025233e-14    2
-3.18909572e+04-1.38313047e+01-4.22291346e-01 3.35894611e-02-2.32937590e-05    3
 8.53864232e-09-1.27783202e-12-2.94428423e+04 2.70882143e+01                   4
N2                      N   2               G    200.00   3500.00 1050.00      1
 2.81166073e+00 1.67067353e-03-6.79997421e-07 1.32881376e-10-1.02767438e-14    2
-8.69811581e+02 6.64838048e+00 3.73100682e+00-1.83159730e-03 4.32324661e-06    3
-3.04378150e-09 7.46071560e-13-1.06287426e+03 2.16821198e+00                   4
O2                      O   2               G    200.00   3500.00  700.00      1
 2.82012408e+00 2.48211357e-03-1.51202094e-06 4.48556199e-10-4.87305665e-14    2
-9.31350152e+02 7.94914552e+00 3.74403921e+00-2.79740146e-03 9.80122556e-06    3
-1.03259643e-08 3.79931246e-12-1.06069827e+03 3.82132646e+00                   4
CO                      C   1O   1          G    200.00   3500.00  960.00      1
 2.79255379e+00 1.87486889e-03-8.59711939e-07 1.91200073e-10-1.67855288e-14    2
-1.41723335e+04 7.41443567e+00 3.75723892e+00-2.14465247e-03 5.42079018e-06    3
-4.17025973e-09 1.11901130e-12-1.43575530e+04 2.79976795e+00                   4
CO2                     C   1O   2          G    200.00   3500.00 1450.00      1
 4.70876459e+00 2.62914723e-03-9.30606600e-07 1.43892961e-10-7.62581846e-15    2
-4.90562638e+04-2.34976404e+00 2.31684348e+00 9.22755029e-03-7.75654080e-06    3
 3.28225351e-09-5.48722465e-13-4.83626067e+04 1.00786234e+01                   4
H2O                     H   2O   1          G    200.00   3500.00 1420.00      1
 2.66777069e+00 3.05768864e-03-9.00442530e-07 1.43361590e-10-1.00857860e-14    2
-2.98875645e+04 6.91191161e+00 4.06061173e+00-8.65807224e-04 3.24409535e-06    3
-1.80243084e-09 3.32483304e-13-3.02831314e+04-2.96150501e-01                   4
END
